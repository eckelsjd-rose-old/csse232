`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:19:45 01/28/2019 
// Design Name: 
// Module Name:    memory_unit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module memory_unit(
	 input clcka,
    input [15:0] a1,
    input [15:0] a2,
    input [15:0] w1,
    input [15:0] w2,
    input w1_ena,
    input w2_ena,
    input r1_ena,
    input r2_ena,
    output [15:0] r1,
    output [15:0] r2,
	 reg
    );

endmodule
